interface adder

logic [6:0]a;
logic [6:0]b;
logic [6:0]c;

endinterface:adder
